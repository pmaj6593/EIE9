`timescale 1 ps / 1 ps
module kernal33_tb(); 

	reg[47:0] im1, im2, im3, k1, k2, k3;
	wire[31:0] result;
	
	kernal33 multi(.im1(im1), .im2(im2), .im3(im3), .k1(k1), .k2(k2), .k3(k3), .result(result));
	
	initial begin
		im1 = 48'b000000000000000100000000000000010000000000000001;
		im2 = 48'b000000000000000100000000000000010000000000000001;
		im3 = 48'b000000000000000100000000000000010000000000000001;
		k1 = 48'b000000000000000100000000000000010000000000000001;
		k2 = 48'b000000000000000100000000000000010000000000000001;
		k3 = 48'b000000000000000100000000000000010000000000000001;
	end

	

endmodule 